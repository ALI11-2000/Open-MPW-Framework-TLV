VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO counter_option1
  CLASS BLOCK ;
  FOREIGN counter_option1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 596.000 8.190 600.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 596.000 242.790 600.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 596.000 266.250 600.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 596.000 289.710 600.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 596.000 313.170 600.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 596.000 336.630 600.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 596.000 360.090 600.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 596.000 383.550 600.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.730 596.000 407.010 600.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 596.000 430.470 600.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 596.000 453.930 600.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 596.000 31.650 600.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 596.000 477.390 600.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.570 596.000 500.850 600.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 596.000 524.310 600.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 596.000 547.770 600.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.950 596.000 571.230 600.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.410 596.000 594.690 600.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.870 596.000 618.150 600.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.330 596.000 641.610 600.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.790 596.000 665.070 600.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 596.000 688.530 600.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 596.000 55.110 600.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 596.000 711.990 600.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.170 596.000 735.450 600.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.630 596.000 758.910 600.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.090 596.000 782.370 600.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.550 596.000 805.830 600.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.010 596.000 829.290 600.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.470 596.000 852.750 600.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.930 596.000 876.210 600.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 596.000 78.570 600.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 596.000 102.030 600.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 596.000 125.490 600.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 596.000 148.950 600.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 596.000 172.410 600.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 596.000 195.870 600.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 596.000 219.330 600.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 596.000 16.010 600.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 596.000 250.610 600.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 596.000 274.070 600.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 596.000 297.530 600.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 596.000 320.990 600.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 596.000 344.450 600.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.630 596.000 367.910 600.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 596.000 391.370 600.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 596.000 414.830 600.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 596.000 438.290 600.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 596.000 461.750 600.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 596.000 39.470 600.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 596.000 485.210 600.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 596.000 508.670 600.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.850 596.000 532.130 600.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.310 596.000 555.590 600.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.770 596.000 579.050 600.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 596.000 602.510 600.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.690 596.000 625.970 600.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.150 596.000 649.430 600.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.610 596.000 672.890 600.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.070 596.000 696.350 600.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 596.000 62.930 600.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.530 596.000 719.810 600.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.990 596.000 743.270 600.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 596.000 766.730 600.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.910 596.000 790.190 600.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.370 596.000 813.650 600.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 836.830 596.000 837.110 600.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.290 596.000 860.570 600.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.750 596.000 884.030 600.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 596.000 86.390 600.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 596.000 109.850 600.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 596.000 133.310 600.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 596.000 156.770 600.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 596.000 180.230 600.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 596.000 203.690 600.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 596.000 227.150 600.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 596.000 23.830 600.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 596.000 258.430 600.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 596.000 281.890 600.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 596.000 305.350 600.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 596.000 328.810 600.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 596.000 352.270 600.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 596.000 375.730 600.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 596.000 399.190 600.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.370 596.000 422.650 600.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.830 596.000 446.110 600.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 596.000 469.570 600.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 596.000 47.290 600.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 596.000 493.030 600.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.210 596.000 516.490 600.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.670 596.000 539.950 600.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.130 596.000 563.410 600.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 596.000 586.870 600.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.050 596.000 610.330 600.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.510 596.000 633.790 600.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 596.000 657.250 600.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.430 596.000 680.710 600.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 596.000 704.170 600.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 596.000 70.750 600.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.350 596.000 727.630 600.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.810 596.000 751.090 600.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.270 596.000 774.550 600.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.730 596.000 798.010 600.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 596.000 821.470 600.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.650 596.000 844.930 600.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.110 596.000 868.390 600.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.570 596.000 891.850 600.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 596.000 94.210 600.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 596.000 117.670 600.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 596.000 141.130 600.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 596.000 164.590 600.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 596.000 188.050 600.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 596.000 211.510 600.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 596.000 234.970 600.000 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.690 0.000 786.970 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.070 0.000 788.350 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.450 0.000 789.730 4.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 0.000 257.050 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.770 0.000 671.050 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 0.000 675.190 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.050 0.000 679.330 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.190 0.000 683.470 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.330 0.000 687.610 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.470 0.000 691.750 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.750 0.000 700.030 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 0.000 704.170 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.030 0.000 708.310 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 0.000 298.450 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.170 0.000 712.450 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.310 0.000 716.590 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.450 0.000 720.730 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 0.000 724.870 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.730 0.000 729.010 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.870 0.000 733.150 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 0.000 737.290 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.150 0.000 741.430 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.290 0.000 745.570 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.430 0.000 749.710 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 0.000 302.590 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 0.000 753.850 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.710 0.000 757.990 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.850 0.000 762.130 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 0.000 766.270 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.130 0.000 770.410 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.270 0.000 774.550 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.410 0.000 778.690 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 0.000 782.830 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 0.000 306.730 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 0.000 310.870 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 0.000 315.010 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 0.000 327.430 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 0.000 331.570 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 0.000 335.710 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 0.000 339.850 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 0.000 343.990 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 0.000 352.270 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 0.000 356.410 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 0.000 360.550 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.550 0.000 368.830 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 0.000 372.970 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 0.000 265.330 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 0.000 381.250 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 0.000 385.390 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 0.000 393.670 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.530 0.000 397.810 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 0.000 401.950 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.950 0.000 410.230 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 0.000 414.370 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 0.000 418.510 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.370 0.000 422.650 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.510 0.000 426.790 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 0.000 430.930 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 0.000 439.210 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 0.000 443.350 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 0.000 447.490 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.350 0.000 451.630 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.490 0.000 455.770 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.630 0.000 459.910 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 0.000 468.190 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.050 0.000 472.330 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 0.000 476.470 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.330 0.000 480.610 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.470 0.000 484.750 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 0.000 488.890 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 0.000 497.170 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.030 0.000 501.310 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 0.000 277.750 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.170 0.000 505.450 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.310 0.000 509.590 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.450 0.000 513.730 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 0.000 517.870 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 0.000 522.010 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.870 0.000 526.150 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 0.000 530.290 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.150 0.000 534.430 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.290 0.000 538.570 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 0.000 542.710 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 0.000 281.890 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.570 0.000 546.850 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 0.000 550.990 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.850 0.000 555.130 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.990 0.000 559.270 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.130 0.000 563.410 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.270 0.000 567.550 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 0.000 571.690 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.550 0.000 575.830 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 0.000 579.970 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.830 0.000 584.110 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 0.000 286.030 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.970 0.000 588.250 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.110 0.000 592.390 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.250 0.000 596.530 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.390 0.000 600.670 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 0.000 604.810 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 0.000 608.950 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 0.000 613.090 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.950 0.000 617.230 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.090 0.000 621.370 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.230 0.000 625.510 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.370 0.000 629.650 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.510 0.000 633.790 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 0.000 637.930 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.790 0.000 642.070 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.930 0.000 646.210 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.070 0.000 650.350 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.210 0.000 654.490 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.350 0.000 658.630 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.490 0.000 662.770 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 0.000 666.910 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 0.000 294.310 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 0.000 258.430 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.150 0.000 672.430 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 0.000 676.570 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.430 0.000 680.710 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.570 0.000 684.850 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.710 0.000 688.990 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.850 0.000 693.130 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.990 0.000 697.270 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.130 0.000 701.410 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 0.000 705.550 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.410 0.000 709.690 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.550 0.000 713.830 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.690 0.000 717.970 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.830 0.000 722.110 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.970 0.000 726.250 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.110 0.000 730.390 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 0.000 734.530 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.390 0.000 738.670 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.530 0.000 742.810 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.670 0.000 746.950 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.810 0.000 751.090 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 0.000 303.970 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.950 0.000 755.230 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.090 0.000 759.370 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 0.000 763.510 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 0.000 767.650 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.510 0.000 771.790 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 0.000 775.930 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.790 0.000 780.070 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.930 0.000 784.210 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 0.000 308.110 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 0.000 312.250 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 0.000 320.530 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 0.000 324.670 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 0.000 332.950 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 0.000 337.090 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 0.000 341.230 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 0.000 345.370 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 0.000 349.510 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.370 0.000 353.650 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 0.000 361.930 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 0.000 366.070 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 0.000 370.210 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.070 0.000 374.350 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 0.000 266.710 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 0.000 382.630 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 0.000 390.910 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 0.000 395.050 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 0.000 399.190 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 0.000 403.330 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 0.000 407.470 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 0.000 411.610 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 0.000 415.750 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.610 0.000 419.890 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.750 0.000 424.030 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 0.000 428.170 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 0.000 432.310 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 0.000 436.450 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 0.000 440.590 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.590 0.000 448.870 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.730 0.000 453.010 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.870 0.000 457.150 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 0.000 461.290 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.150 0.000 465.430 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 0.000 469.570 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.570 0.000 477.850 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 0.000 481.990 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 0.000 486.130 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.990 0.000 490.270 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.130 0.000 494.410 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.270 0.000 498.550 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 0.000 279.130 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.550 0.000 506.830 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 0.000 510.970 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 0.000 515.110 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.970 0.000 519.250 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.110 0.000 523.390 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.250 0.000 527.530 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 0.000 535.810 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.670 0.000 539.950 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 0.000 544.090 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 0.000 283.270 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 0.000 548.230 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 0.000 552.370 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 0.000 556.510 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 0.000 564.790 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.650 0.000 568.930 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.790 0.000 573.070 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.930 0.000 577.210 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 0.000 581.350 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 0.000 585.490 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 0.000 287.410 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.490 0.000 593.770 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 0.000 597.910 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.770 0.000 602.050 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.910 0.000 606.190 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.050 0.000 610.330 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.190 0.000 614.470 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 0.000 618.610 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.470 0.000 622.750 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.610 0.000 626.890 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 0.000 291.550 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.750 0.000 631.030 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.890 0.000 635.170 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.030 0.000 639.310 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.170 0.000 643.450 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 0.000 647.590 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.450 0.000 651.730 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.590 0.000 655.870 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.730 0.000 660.010 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.870 0.000 664.150 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.010 0.000 668.290 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.530 0.000 673.810 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.670 0.000 677.950 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.810 0.000 682.090 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 0.000 686.230 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.090 0.000 690.370 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 0.000 694.510 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.370 0.000 698.650 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 0.000 702.790 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.650 0.000 706.930 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.790 0.000 711.070 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 0.000 301.210 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.070 0.000 719.350 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.210 0.000 723.490 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.350 0.000 727.630 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.490 0.000 731.770 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.630 0.000 735.910 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.770 0.000 740.050 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 0.000 744.190 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.050 0.000 748.330 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.190 0.000 752.470 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 0.000 305.350 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.330 0.000 756.610 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.470 0.000 760.750 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.610 0.000 764.890 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.750 0.000 769.030 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 0.000 773.170 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.030 0.000 777.310 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.170 0.000 781.450 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.310 0.000 785.590 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 0.000 313.630 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 0.000 321.910 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 0.000 330.190 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 0.000 346.750 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 0.000 350.890 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 0.000 355.030 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 0.000 359.170 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.030 0.000 363.310 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 0.000 371.590 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 0.000 375.730 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 0.000 379.870 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.730 0.000 384.010 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 0.000 388.150 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 0.000 400.570 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.430 0.000 404.710 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.570 0.000 408.850 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 0.000 412.990 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.850 0.000 417.130 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 0.000 421.270 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 0.000 272.230 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 0.000 429.550 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.410 0.000 433.690 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 0.000 437.830 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 0.000 441.970 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.830 0.000 446.110 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 0.000 450.250 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 0.000 458.530 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 0.000 462.670 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.530 0.000 466.810 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.670 0.000 470.950 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.810 0.000 475.090 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 0.000 487.510 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 0.000 491.650 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 0.000 495.790 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 0.000 499.930 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.790 0.000 504.070 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.930 0.000 508.210 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.210 0.000 516.490 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.350 0.000 520.630 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 0.000 524.770 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.630 0.000 528.910 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.770 0.000 533.050 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.910 0.000 537.190 4.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 0.000 541.330 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.190 0.000 545.470 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.330 0.000 549.610 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 0.000 553.750 4.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.610 0.000 557.890 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.750 0.000 562.030 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.890 0.000 566.170 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 0.000 570.310 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.170 0.000 574.450 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 0.000 578.590 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.450 0.000 582.730 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 0.000 586.870 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.730 0.000 591.010 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.870 0.000 595.150 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.150 0.000 603.430 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.290 0.000 607.570 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.430 0.000 611.710 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.570 0.000 615.850 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.710 0.000 619.990 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 0.000 624.130 4.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 0.000 628.270 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130 0.000 632.410 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.270 0.000 636.550 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.410 0.000 640.690 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.550 0.000 644.830 4.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.690 0.000 648.970 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.830 0.000 653.110 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 0.000 657.250 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.110 0.000 661.390 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.250 0.000 665.530 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.390 0.000 669.670 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END la_oenb[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 587.760 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 0.000 170.110 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 0.000 186.670 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 0.000 211.510 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 0.000 219.790 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 0.000 223.930 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 0.000 244.630 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.770 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 0.000 252.910 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 0.000 153.550 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 0.000 167.350 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 0.000 196.330 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 0.000 204.610 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 0.000 217.030 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 0.000 229.450 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 0.000 233.590 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 0.000 181.150 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.430 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 0.000 239.110 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 0.000 148.030 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 0.000 128.710 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER nwell ;
        RECT 5.330 583.385 894.430 586.215 ;
        RECT 5.330 577.945 894.430 580.775 ;
        RECT 5.330 572.505 894.430 575.335 ;
        RECT 5.330 567.065 894.430 569.895 ;
        RECT 5.330 561.625 894.430 564.455 ;
        RECT 5.330 556.185 894.430 559.015 ;
        RECT 5.330 550.745 894.430 553.575 ;
        RECT 5.330 545.305 894.430 548.135 ;
        RECT 5.330 539.865 894.430 542.695 ;
        RECT 5.330 534.425 894.430 537.255 ;
        RECT 5.330 528.985 894.430 531.815 ;
        RECT 5.330 523.545 894.430 526.375 ;
        RECT 5.330 518.105 894.430 520.935 ;
        RECT 5.330 512.665 894.430 515.495 ;
        RECT 5.330 507.225 894.430 510.055 ;
        RECT 5.330 501.785 894.430 504.615 ;
        RECT 5.330 496.345 894.430 499.175 ;
        RECT 5.330 490.905 894.430 493.735 ;
        RECT 5.330 485.465 894.430 488.295 ;
        RECT 5.330 480.025 894.430 482.855 ;
        RECT 5.330 474.585 894.430 477.415 ;
        RECT 5.330 469.145 894.430 471.975 ;
        RECT 5.330 463.705 894.430 466.535 ;
        RECT 5.330 458.265 894.430 461.095 ;
        RECT 5.330 452.825 894.430 455.655 ;
        RECT 5.330 447.385 894.430 450.215 ;
        RECT 5.330 441.945 894.430 444.775 ;
        RECT 5.330 436.505 894.430 439.335 ;
        RECT 5.330 431.065 894.430 433.895 ;
        RECT 5.330 425.625 894.430 428.455 ;
        RECT 5.330 420.185 894.430 423.015 ;
        RECT 5.330 414.745 894.430 417.575 ;
        RECT 5.330 409.305 894.430 412.135 ;
        RECT 5.330 403.865 894.430 406.695 ;
        RECT 5.330 398.425 894.430 401.255 ;
        RECT 5.330 392.985 894.430 395.815 ;
        RECT 5.330 387.545 894.430 390.375 ;
        RECT 5.330 382.105 894.430 384.935 ;
        RECT 5.330 376.665 894.430 379.495 ;
        RECT 5.330 371.225 894.430 374.055 ;
        RECT 5.330 365.785 894.430 368.615 ;
        RECT 5.330 360.345 894.430 363.175 ;
        RECT 5.330 354.905 894.430 357.735 ;
        RECT 5.330 349.465 894.430 352.295 ;
        RECT 5.330 344.025 894.430 346.855 ;
        RECT 5.330 338.585 894.430 341.415 ;
        RECT 5.330 333.145 894.430 335.975 ;
        RECT 5.330 327.705 894.430 330.535 ;
        RECT 5.330 322.265 894.430 325.095 ;
        RECT 5.330 316.825 894.430 319.655 ;
        RECT 5.330 311.385 894.430 314.215 ;
        RECT 5.330 305.945 894.430 308.775 ;
        RECT 5.330 300.505 894.430 303.335 ;
        RECT 5.330 295.065 894.430 297.895 ;
        RECT 5.330 289.625 894.430 292.455 ;
        RECT 5.330 284.185 894.430 287.015 ;
        RECT 5.330 278.745 894.430 281.575 ;
        RECT 5.330 273.305 894.430 276.135 ;
        RECT 5.330 267.865 894.430 270.695 ;
        RECT 5.330 262.425 894.430 265.255 ;
        RECT 5.330 256.985 894.430 259.815 ;
        RECT 5.330 251.545 894.430 254.375 ;
        RECT 5.330 246.105 894.430 248.935 ;
        RECT 5.330 240.665 894.430 243.495 ;
        RECT 5.330 235.225 894.430 238.055 ;
        RECT 5.330 229.785 894.430 232.615 ;
        RECT 5.330 224.345 894.430 227.175 ;
        RECT 5.330 218.905 894.430 221.735 ;
        RECT 5.330 213.465 894.430 216.295 ;
        RECT 5.330 208.025 894.430 210.855 ;
        RECT 5.330 202.585 894.430 205.415 ;
        RECT 5.330 197.145 894.430 199.975 ;
        RECT 5.330 191.705 894.430 194.535 ;
        RECT 5.330 186.265 894.430 189.095 ;
        RECT 5.330 180.825 894.430 183.655 ;
        RECT 5.330 175.385 894.430 178.215 ;
        RECT 5.330 169.945 894.430 172.775 ;
        RECT 5.330 164.505 894.430 167.335 ;
        RECT 5.330 159.065 894.430 161.895 ;
        RECT 5.330 153.625 894.430 156.455 ;
        RECT 5.330 148.185 894.430 151.015 ;
        RECT 5.330 142.745 894.430 145.575 ;
        RECT 5.330 137.305 894.430 140.135 ;
        RECT 5.330 131.865 894.430 134.695 ;
        RECT 5.330 126.425 894.430 129.255 ;
        RECT 5.330 120.985 894.430 123.815 ;
        RECT 5.330 115.545 894.430 118.375 ;
        RECT 5.330 110.105 894.430 112.935 ;
        RECT 5.330 104.665 894.430 107.495 ;
        RECT 5.330 99.225 894.430 102.055 ;
        RECT 5.330 93.785 894.430 96.615 ;
        RECT 5.330 88.345 894.430 91.175 ;
        RECT 5.330 82.905 894.430 85.735 ;
        RECT 5.330 77.465 894.430 80.295 ;
        RECT 5.330 72.025 894.430 74.855 ;
        RECT 5.330 66.585 894.430 69.415 ;
        RECT 5.330 61.145 894.430 63.975 ;
        RECT 5.330 55.705 894.430 58.535 ;
        RECT 5.330 50.265 894.430 53.095 ;
        RECT 5.330 44.825 894.430 47.655 ;
        RECT 5.330 39.385 894.430 42.215 ;
        RECT 5.330 33.945 894.430 36.775 ;
        RECT 5.330 28.505 894.430 31.335 ;
        RECT 5.330 23.065 894.430 25.895 ;
        RECT 5.330 17.625 894.430 20.455 ;
        RECT 5.330 12.185 894.430 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 894.240 587.605 ;
      LAYER met1 ;
        RECT 5.520 8.880 894.240 587.760 ;
      LAYER met2 ;
        RECT 16.290 595.720 23.270 596.770 ;
        RECT 24.110 595.720 31.090 596.770 ;
        RECT 31.930 595.720 38.910 596.770 ;
        RECT 39.750 595.720 46.730 596.770 ;
        RECT 47.570 595.720 54.550 596.770 ;
        RECT 55.390 595.720 62.370 596.770 ;
        RECT 63.210 595.720 70.190 596.770 ;
        RECT 71.030 595.720 78.010 596.770 ;
        RECT 78.850 595.720 85.830 596.770 ;
        RECT 86.670 595.720 93.650 596.770 ;
        RECT 94.490 595.720 101.470 596.770 ;
        RECT 102.310 595.720 109.290 596.770 ;
        RECT 110.130 595.720 117.110 596.770 ;
        RECT 117.950 595.720 124.930 596.770 ;
        RECT 125.770 595.720 132.750 596.770 ;
        RECT 133.590 595.720 140.570 596.770 ;
        RECT 141.410 595.720 148.390 596.770 ;
        RECT 149.230 595.720 156.210 596.770 ;
        RECT 157.050 595.720 164.030 596.770 ;
        RECT 164.870 595.720 171.850 596.770 ;
        RECT 172.690 595.720 179.670 596.770 ;
        RECT 180.510 595.720 187.490 596.770 ;
        RECT 188.330 595.720 195.310 596.770 ;
        RECT 196.150 595.720 203.130 596.770 ;
        RECT 203.970 595.720 210.950 596.770 ;
        RECT 211.790 595.720 218.770 596.770 ;
        RECT 219.610 595.720 226.590 596.770 ;
        RECT 227.430 595.720 234.410 596.770 ;
        RECT 235.250 595.720 242.230 596.770 ;
        RECT 243.070 595.720 250.050 596.770 ;
        RECT 250.890 595.720 257.870 596.770 ;
        RECT 258.710 595.720 265.690 596.770 ;
        RECT 266.530 595.720 273.510 596.770 ;
        RECT 274.350 595.720 281.330 596.770 ;
        RECT 282.170 595.720 289.150 596.770 ;
        RECT 289.990 595.720 296.970 596.770 ;
        RECT 297.810 595.720 304.790 596.770 ;
        RECT 305.630 595.720 312.610 596.770 ;
        RECT 313.450 595.720 320.430 596.770 ;
        RECT 321.270 595.720 328.250 596.770 ;
        RECT 329.090 595.720 336.070 596.770 ;
        RECT 336.910 595.720 343.890 596.770 ;
        RECT 344.730 595.720 351.710 596.770 ;
        RECT 352.550 595.720 359.530 596.770 ;
        RECT 360.370 595.720 367.350 596.770 ;
        RECT 368.190 595.720 375.170 596.770 ;
        RECT 376.010 595.720 382.990 596.770 ;
        RECT 383.830 595.720 390.810 596.770 ;
        RECT 391.650 595.720 398.630 596.770 ;
        RECT 399.470 595.720 406.450 596.770 ;
        RECT 407.290 595.720 414.270 596.770 ;
        RECT 415.110 595.720 422.090 596.770 ;
        RECT 422.930 595.720 429.910 596.770 ;
        RECT 430.750 595.720 437.730 596.770 ;
        RECT 438.570 595.720 445.550 596.770 ;
        RECT 446.390 595.720 453.370 596.770 ;
        RECT 454.210 595.720 461.190 596.770 ;
        RECT 462.030 595.720 469.010 596.770 ;
        RECT 469.850 595.720 476.830 596.770 ;
        RECT 477.670 595.720 484.650 596.770 ;
        RECT 485.490 595.720 492.470 596.770 ;
        RECT 493.310 595.720 500.290 596.770 ;
        RECT 501.130 595.720 508.110 596.770 ;
        RECT 508.950 595.720 515.930 596.770 ;
        RECT 516.770 595.720 523.750 596.770 ;
        RECT 524.590 595.720 531.570 596.770 ;
        RECT 532.410 595.720 539.390 596.770 ;
        RECT 540.230 595.720 547.210 596.770 ;
        RECT 548.050 595.720 555.030 596.770 ;
        RECT 555.870 595.720 562.850 596.770 ;
        RECT 563.690 595.720 570.670 596.770 ;
        RECT 571.510 595.720 578.490 596.770 ;
        RECT 579.330 595.720 586.310 596.770 ;
        RECT 587.150 595.720 594.130 596.770 ;
        RECT 594.970 595.720 601.950 596.770 ;
        RECT 602.790 595.720 609.770 596.770 ;
        RECT 610.610 595.720 617.590 596.770 ;
        RECT 618.430 595.720 625.410 596.770 ;
        RECT 626.250 595.720 633.230 596.770 ;
        RECT 634.070 595.720 641.050 596.770 ;
        RECT 641.890 595.720 648.870 596.770 ;
        RECT 649.710 595.720 656.690 596.770 ;
        RECT 657.530 595.720 664.510 596.770 ;
        RECT 665.350 595.720 672.330 596.770 ;
        RECT 673.170 595.720 680.150 596.770 ;
        RECT 680.990 595.720 687.970 596.770 ;
        RECT 688.810 595.720 695.790 596.770 ;
        RECT 696.630 595.720 703.610 596.770 ;
        RECT 704.450 595.720 711.430 596.770 ;
        RECT 712.270 595.720 719.250 596.770 ;
        RECT 720.090 595.720 727.070 596.770 ;
        RECT 727.910 595.720 734.890 596.770 ;
        RECT 735.730 595.720 742.710 596.770 ;
        RECT 743.550 595.720 750.530 596.770 ;
        RECT 751.370 595.720 758.350 596.770 ;
        RECT 759.190 595.720 766.170 596.770 ;
        RECT 767.010 595.720 773.990 596.770 ;
        RECT 774.830 595.720 781.810 596.770 ;
        RECT 782.650 595.720 789.630 596.770 ;
        RECT 790.470 595.720 797.450 596.770 ;
        RECT 798.290 595.720 805.270 596.770 ;
        RECT 806.110 595.720 813.090 596.770 ;
        RECT 813.930 595.720 820.910 596.770 ;
        RECT 821.750 595.720 828.730 596.770 ;
        RECT 829.570 595.720 836.550 596.770 ;
        RECT 837.390 595.720 844.370 596.770 ;
        RECT 845.210 595.720 852.190 596.770 ;
        RECT 853.030 595.720 860.010 596.770 ;
        RECT 860.850 595.720 867.830 596.770 ;
        RECT 868.670 595.720 875.650 596.770 ;
        RECT 876.490 595.720 883.470 596.770 ;
        RECT 884.310 595.720 891.290 596.770 ;
        RECT 15.740 4.280 891.570 595.720 ;
        RECT 15.740 3.670 110.210 4.280 ;
        RECT 111.050 3.670 111.590 4.280 ;
        RECT 112.430 3.670 112.970 4.280 ;
        RECT 113.810 3.670 114.350 4.280 ;
        RECT 115.190 3.670 115.730 4.280 ;
        RECT 116.570 3.670 117.110 4.280 ;
        RECT 117.950 3.670 118.490 4.280 ;
        RECT 119.330 3.670 119.870 4.280 ;
        RECT 120.710 3.670 121.250 4.280 ;
        RECT 122.090 3.670 122.630 4.280 ;
        RECT 123.470 3.670 124.010 4.280 ;
        RECT 124.850 3.670 125.390 4.280 ;
        RECT 126.230 3.670 126.770 4.280 ;
        RECT 127.610 3.670 128.150 4.280 ;
        RECT 128.990 3.670 129.530 4.280 ;
        RECT 130.370 3.670 130.910 4.280 ;
        RECT 131.750 3.670 132.290 4.280 ;
        RECT 133.130 3.670 133.670 4.280 ;
        RECT 134.510 3.670 135.050 4.280 ;
        RECT 135.890 3.670 136.430 4.280 ;
        RECT 137.270 3.670 137.810 4.280 ;
        RECT 138.650 3.670 139.190 4.280 ;
        RECT 140.030 3.670 140.570 4.280 ;
        RECT 141.410 3.670 141.950 4.280 ;
        RECT 142.790 3.670 143.330 4.280 ;
        RECT 144.170 3.670 144.710 4.280 ;
        RECT 145.550 3.670 146.090 4.280 ;
        RECT 146.930 3.670 147.470 4.280 ;
        RECT 148.310 3.670 148.850 4.280 ;
        RECT 149.690 3.670 150.230 4.280 ;
        RECT 151.070 3.670 151.610 4.280 ;
        RECT 152.450 3.670 152.990 4.280 ;
        RECT 153.830 3.670 154.370 4.280 ;
        RECT 155.210 3.670 155.750 4.280 ;
        RECT 156.590 3.670 157.130 4.280 ;
        RECT 157.970 3.670 158.510 4.280 ;
        RECT 159.350 3.670 159.890 4.280 ;
        RECT 160.730 3.670 161.270 4.280 ;
        RECT 162.110 3.670 162.650 4.280 ;
        RECT 163.490 3.670 164.030 4.280 ;
        RECT 164.870 3.670 165.410 4.280 ;
        RECT 166.250 3.670 166.790 4.280 ;
        RECT 167.630 3.670 168.170 4.280 ;
        RECT 169.010 3.670 169.550 4.280 ;
        RECT 170.390 3.670 170.930 4.280 ;
        RECT 171.770 3.670 172.310 4.280 ;
        RECT 173.150 3.670 173.690 4.280 ;
        RECT 174.530 3.670 175.070 4.280 ;
        RECT 175.910 3.670 176.450 4.280 ;
        RECT 177.290 3.670 177.830 4.280 ;
        RECT 178.670 3.670 179.210 4.280 ;
        RECT 180.050 3.670 180.590 4.280 ;
        RECT 181.430 3.670 181.970 4.280 ;
        RECT 182.810 3.670 183.350 4.280 ;
        RECT 184.190 3.670 184.730 4.280 ;
        RECT 185.570 3.670 186.110 4.280 ;
        RECT 186.950 3.670 187.490 4.280 ;
        RECT 188.330 3.670 188.870 4.280 ;
        RECT 189.710 3.670 190.250 4.280 ;
        RECT 191.090 3.670 191.630 4.280 ;
        RECT 192.470 3.670 193.010 4.280 ;
        RECT 193.850 3.670 194.390 4.280 ;
        RECT 195.230 3.670 195.770 4.280 ;
        RECT 196.610 3.670 197.150 4.280 ;
        RECT 197.990 3.670 198.530 4.280 ;
        RECT 199.370 3.670 199.910 4.280 ;
        RECT 200.750 3.670 201.290 4.280 ;
        RECT 202.130 3.670 202.670 4.280 ;
        RECT 203.510 3.670 204.050 4.280 ;
        RECT 204.890 3.670 205.430 4.280 ;
        RECT 206.270 3.670 206.810 4.280 ;
        RECT 207.650 3.670 208.190 4.280 ;
        RECT 209.030 3.670 209.570 4.280 ;
        RECT 210.410 3.670 210.950 4.280 ;
        RECT 211.790 3.670 212.330 4.280 ;
        RECT 213.170 3.670 213.710 4.280 ;
        RECT 214.550 3.670 215.090 4.280 ;
        RECT 215.930 3.670 216.470 4.280 ;
        RECT 217.310 3.670 217.850 4.280 ;
        RECT 218.690 3.670 219.230 4.280 ;
        RECT 220.070 3.670 220.610 4.280 ;
        RECT 221.450 3.670 221.990 4.280 ;
        RECT 222.830 3.670 223.370 4.280 ;
        RECT 224.210 3.670 224.750 4.280 ;
        RECT 225.590 3.670 226.130 4.280 ;
        RECT 226.970 3.670 227.510 4.280 ;
        RECT 228.350 3.670 228.890 4.280 ;
        RECT 229.730 3.670 230.270 4.280 ;
        RECT 231.110 3.670 231.650 4.280 ;
        RECT 232.490 3.670 233.030 4.280 ;
        RECT 233.870 3.670 234.410 4.280 ;
        RECT 235.250 3.670 235.790 4.280 ;
        RECT 236.630 3.670 237.170 4.280 ;
        RECT 238.010 3.670 238.550 4.280 ;
        RECT 239.390 3.670 239.930 4.280 ;
        RECT 240.770 3.670 241.310 4.280 ;
        RECT 242.150 3.670 242.690 4.280 ;
        RECT 243.530 3.670 244.070 4.280 ;
        RECT 244.910 3.670 245.450 4.280 ;
        RECT 246.290 3.670 246.830 4.280 ;
        RECT 247.670 3.670 248.210 4.280 ;
        RECT 249.050 3.670 249.590 4.280 ;
        RECT 250.430 3.670 250.970 4.280 ;
        RECT 251.810 3.670 252.350 4.280 ;
        RECT 253.190 3.670 253.730 4.280 ;
        RECT 254.570 3.670 255.110 4.280 ;
        RECT 255.950 3.670 256.490 4.280 ;
        RECT 257.330 3.670 257.870 4.280 ;
        RECT 258.710 3.670 259.250 4.280 ;
        RECT 260.090 3.670 260.630 4.280 ;
        RECT 261.470 3.670 262.010 4.280 ;
        RECT 262.850 3.670 263.390 4.280 ;
        RECT 264.230 3.670 264.770 4.280 ;
        RECT 265.610 3.670 266.150 4.280 ;
        RECT 266.990 3.670 267.530 4.280 ;
        RECT 268.370 3.670 268.910 4.280 ;
        RECT 269.750 3.670 270.290 4.280 ;
        RECT 271.130 3.670 271.670 4.280 ;
        RECT 272.510 3.670 273.050 4.280 ;
        RECT 273.890 3.670 274.430 4.280 ;
        RECT 275.270 3.670 275.810 4.280 ;
        RECT 276.650 3.670 277.190 4.280 ;
        RECT 278.030 3.670 278.570 4.280 ;
        RECT 279.410 3.670 279.950 4.280 ;
        RECT 280.790 3.670 281.330 4.280 ;
        RECT 282.170 3.670 282.710 4.280 ;
        RECT 283.550 3.670 284.090 4.280 ;
        RECT 284.930 3.670 285.470 4.280 ;
        RECT 286.310 3.670 286.850 4.280 ;
        RECT 287.690 3.670 288.230 4.280 ;
        RECT 289.070 3.670 289.610 4.280 ;
        RECT 290.450 3.670 290.990 4.280 ;
        RECT 291.830 3.670 292.370 4.280 ;
        RECT 293.210 3.670 293.750 4.280 ;
        RECT 294.590 3.670 295.130 4.280 ;
        RECT 295.970 3.670 296.510 4.280 ;
        RECT 297.350 3.670 297.890 4.280 ;
        RECT 298.730 3.670 299.270 4.280 ;
        RECT 300.110 3.670 300.650 4.280 ;
        RECT 301.490 3.670 302.030 4.280 ;
        RECT 302.870 3.670 303.410 4.280 ;
        RECT 304.250 3.670 304.790 4.280 ;
        RECT 305.630 3.670 306.170 4.280 ;
        RECT 307.010 3.670 307.550 4.280 ;
        RECT 308.390 3.670 308.930 4.280 ;
        RECT 309.770 3.670 310.310 4.280 ;
        RECT 311.150 3.670 311.690 4.280 ;
        RECT 312.530 3.670 313.070 4.280 ;
        RECT 313.910 3.670 314.450 4.280 ;
        RECT 315.290 3.670 315.830 4.280 ;
        RECT 316.670 3.670 317.210 4.280 ;
        RECT 318.050 3.670 318.590 4.280 ;
        RECT 319.430 3.670 319.970 4.280 ;
        RECT 320.810 3.670 321.350 4.280 ;
        RECT 322.190 3.670 322.730 4.280 ;
        RECT 323.570 3.670 324.110 4.280 ;
        RECT 324.950 3.670 325.490 4.280 ;
        RECT 326.330 3.670 326.870 4.280 ;
        RECT 327.710 3.670 328.250 4.280 ;
        RECT 329.090 3.670 329.630 4.280 ;
        RECT 330.470 3.670 331.010 4.280 ;
        RECT 331.850 3.670 332.390 4.280 ;
        RECT 333.230 3.670 333.770 4.280 ;
        RECT 334.610 3.670 335.150 4.280 ;
        RECT 335.990 3.670 336.530 4.280 ;
        RECT 337.370 3.670 337.910 4.280 ;
        RECT 338.750 3.670 339.290 4.280 ;
        RECT 340.130 3.670 340.670 4.280 ;
        RECT 341.510 3.670 342.050 4.280 ;
        RECT 342.890 3.670 343.430 4.280 ;
        RECT 344.270 3.670 344.810 4.280 ;
        RECT 345.650 3.670 346.190 4.280 ;
        RECT 347.030 3.670 347.570 4.280 ;
        RECT 348.410 3.670 348.950 4.280 ;
        RECT 349.790 3.670 350.330 4.280 ;
        RECT 351.170 3.670 351.710 4.280 ;
        RECT 352.550 3.670 353.090 4.280 ;
        RECT 353.930 3.670 354.470 4.280 ;
        RECT 355.310 3.670 355.850 4.280 ;
        RECT 356.690 3.670 357.230 4.280 ;
        RECT 358.070 3.670 358.610 4.280 ;
        RECT 359.450 3.670 359.990 4.280 ;
        RECT 360.830 3.670 361.370 4.280 ;
        RECT 362.210 3.670 362.750 4.280 ;
        RECT 363.590 3.670 364.130 4.280 ;
        RECT 364.970 3.670 365.510 4.280 ;
        RECT 366.350 3.670 366.890 4.280 ;
        RECT 367.730 3.670 368.270 4.280 ;
        RECT 369.110 3.670 369.650 4.280 ;
        RECT 370.490 3.670 371.030 4.280 ;
        RECT 371.870 3.670 372.410 4.280 ;
        RECT 373.250 3.670 373.790 4.280 ;
        RECT 374.630 3.670 375.170 4.280 ;
        RECT 376.010 3.670 376.550 4.280 ;
        RECT 377.390 3.670 377.930 4.280 ;
        RECT 378.770 3.670 379.310 4.280 ;
        RECT 380.150 3.670 380.690 4.280 ;
        RECT 381.530 3.670 382.070 4.280 ;
        RECT 382.910 3.670 383.450 4.280 ;
        RECT 384.290 3.670 384.830 4.280 ;
        RECT 385.670 3.670 386.210 4.280 ;
        RECT 387.050 3.670 387.590 4.280 ;
        RECT 388.430 3.670 388.970 4.280 ;
        RECT 389.810 3.670 390.350 4.280 ;
        RECT 391.190 3.670 391.730 4.280 ;
        RECT 392.570 3.670 393.110 4.280 ;
        RECT 393.950 3.670 394.490 4.280 ;
        RECT 395.330 3.670 395.870 4.280 ;
        RECT 396.710 3.670 397.250 4.280 ;
        RECT 398.090 3.670 398.630 4.280 ;
        RECT 399.470 3.670 400.010 4.280 ;
        RECT 400.850 3.670 401.390 4.280 ;
        RECT 402.230 3.670 402.770 4.280 ;
        RECT 403.610 3.670 404.150 4.280 ;
        RECT 404.990 3.670 405.530 4.280 ;
        RECT 406.370 3.670 406.910 4.280 ;
        RECT 407.750 3.670 408.290 4.280 ;
        RECT 409.130 3.670 409.670 4.280 ;
        RECT 410.510 3.670 411.050 4.280 ;
        RECT 411.890 3.670 412.430 4.280 ;
        RECT 413.270 3.670 413.810 4.280 ;
        RECT 414.650 3.670 415.190 4.280 ;
        RECT 416.030 3.670 416.570 4.280 ;
        RECT 417.410 3.670 417.950 4.280 ;
        RECT 418.790 3.670 419.330 4.280 ;
        RECT 420.170 3.670 420.710 4.280 ;
        RECT 421.550 3.670 422.090 4.280 ;
        RECT 422.930 3.670 423.470 4.280 ;
        RECT 424.310 3.670 424.850 4.280 ;
        RECT 425.690 3.670 426.230 4.280 ;
        RECT 427.070 3.670 427.610 4.280 ;
        RECT 428.450 3.670 428.990 4.280 ;
        RECT 429.830 3.670 430.370 4.280 ;
        RECT 431.210 3.670 431.750 4.280 ;
        RECT 432.590 3.670 433.130 4.280 ;
        RECT 433.970 3.670 434.510 4.280 ;
        RECT 435.350 3.670 435.890 4.280 ;
        RECT 436.730 3.670 437.270 4.280 ;
        RECT 438.110 3.670 438.650 4.280 ;
        RECT 439.490 3.670 440.030 4.280 ;
        RECT 440.870 3.670 441.410 4.280 ;
        RECT 442.250 3.670 442.790 4.280 ;
        RECT 443.630 3.670 444.170 4.280 ;
        RECT 445.010 3.670 445.550 4.280 ;
        RECT 446.390 3.670 446.930 4.280 ;
        RECT 447.770 3.670 448.310 4.280 ;
        RECT 449.150 3.670 449.690 4.280 ;
        RECT 450.530 3.670 451.070 4.280 ;
        RECT 451.910 3.670 452.450 4.280 ;
        RECT 453.290 3.670 453.830 4.280 ;
        RECT 454.670 3.670 455.210 4.280 ;
        RECT 456.050 3.670 456.590 4.280 ;
        RECT 457.430 3.670 457.970 4.280 ;
        RECT 458.810 3.670 459.350 4.280 ;
        RECT 460.190 3.670 460.730 4.280 ;
        RECT 461.570 3.670 462.110 4.280 ;
        RECT 462.950 3.670 463.490 4.280 ;
        RECT 464.330 3.670 464.870 4.280 ;
        RECT 465.710 3.670 466.250 4.280 ;
        RECT 467.090 3.670 467.630 4.280 ;
        RECT 468.470 3.670 469.010 4.280 ;
        RECT 469.850 3.670 470.390 4.280 ;
        RECT 471.230 3.670 471.770 4.280 ;
        RECT 472.610 3.670 473.150 4.280 ;
        RECT 473.990 3.670 474.530 4.280 ;
        RECT 475.370 3.670 475.910 4.280 ;
        RECT 476.750 3.670 477.290 4.280 ;
        RECT 478.130 3.670 478.670 4.280 ;
        RECT 479.510 3.670 480.050 4.280 ;
        RECT 480.890 3.670 481.430 4.280 ;
        RECT 482.270 3.670 482.810 4.280 ;
        RECT 483.650 3.670 484.190 4.280 ;
        RECT 485.030 3.670 485.570 4.280 ;
        RECT 486.410 3.670 486.950 4.280 ;
        RECT 487.790 3.670 488.330 4.280 ;
        RECT 489.170 3.670 489.710 4.280 ;
        RECT 490.550 3.670 491.090 4.280 ;
        RECT 491.930 3.670 492.470 4.280 ;
        RECT 493.310 3.670 493.850 4.280 ;
        RECT 494.690 3.670 495.230 4.280 ;
        RECT 496.070 3.670 496.610 4.280 ;
        RECT 497.450 3.670 497.990 4.280 ;
        RECT 498.830 3.670 499.370 4.280 ;
        RECT 500.210 3.670 500.750 4.280 ;
        RECT 501.590 3.670 502.130 4.280 ;
        RECT 502.970 3.670 503.510 4.280 ;
        RECT 504.350 3.670 504.890 4.280 ;
        RECT 505.730 3.670 506.270 4.280 ;
        RECT 507.110 3.670 507.650 4.280 ;
        RECT 508.490 3.670 509.030 4.280 ;
        RECT 509.870 3.670 510.410 4.280 ;
        RECT 511.250 3.670 511.790 4.280 ;
        RECT 512.630 3.670 513.170 4.280 ;
        RECT 514.010 3.670 514.550 4.280 ;
        RECT 515.390 3.670 515.930 4.280 ;
        RECT 516.770 3.670 517.310 4.280 ;
        RECT 518.150 3.670 518.690 4.280 ;
        RECT 519.530 3.670 520.070 4.280 ;
        RECT 520.910 3.670 521.450 4.280 ;
        RECT 522.290 3.670 522.830 4.280 ;
        RECT 523.670 3.670 524.210 4.280 ;
        RECT 525.050 3.670 525.590 4.280 ;
        RECT 526.430 3.670 526.970 4.280 ;
        RECT 527.810 3.670 528.350 4.280 ;
        RECT 529.190 3.670 529.730 4.280 ;
        RECT 530.570 3.670 531.110 4.280 ;
        RECT 531.950 3.670 532.490 4.280 ;
        RECT 533.330 3.670 533.870 4.280 ;
        RECT 534.710 3.670 535.250 4.280 ;
        RECT 536.090 3.670 536.630 4.280 ;
        RECT 537.470 3.670 538.010 4.280 ;
        RECT 538.850 3.670 539.390 4.280 ;
        RECT 540.230 3.670 540.770 4.280 ;
        RECT 541.610 3.670 542.150 4.280 ;
        RECT 542.990 3.670 543.530 4.280 ;
        RECT 544.370 3.670 544.910 4.280 ;
        RECT 545.750 3.670 546.290 4.280 ;
        RECT 547.130 3.670 547.670 4.280 ;
        RECT 548.510 3.670 549.050 4.280 ;
        RECT 549.890 3.670 550.430 4.280 ;
        RECT 551.270 3.670 551.810 4.280 ;
        RECT 552.650 3.670 553.190 4.280 ;
        RECT 554.030 3.670 554.570 4.280 ;
        RECT 555.410 3.670 555.950 4.280 ;
        RECT 556.790 3.670 557.330 4.280 ;
        RECT 558.170 3.670 558.710 4.280 ;
        RECT 559.550 3.670 560.090 4.280 ;
        RECT 560.930 3.670 561.470 4.280 ;
        RECT 562.310 3.670 562.850 4.280 ;
        RECT 563.690 3.670 564.230 4.280 ;
        RECT 565.070 3.670 565.610 4.280 ;
        RECT 566.450 3.670 566.990 4.280 ;
        RECT 567.830 3.670 568.370 4.280 ;
        RECT 569.210 3.670 569.750 4.280 ;
        RECT 570.590 3.670 571.130 4.280 ;
        RECT 571.970 3.670 572.510 4.280 ;
        RECT 573.350 3.670 573.890 4.280 ;
        RECT 574.730 3.670 575.270 4.280 ;
        RECT 576.110 3.670 576.650 4.280 ;
        RECT 577.490 3.670 578.030 4.280 ;
        RECT 578.870 3.670 579.410 4.280 ;
        RECT 580.250 3.670 580.790 4.280 ;
        RECT 581.630 3.670 582.170 4.280 ;
        RECT 583.010 3.670 583.550 4.280 ;
        RECT 584.390 3.670 584.930 4.280 ;
        RECT 585.770 3.670 586.310 4.280 ;
        RECT 587.150 3.670 587.690 4.280 ;
        RECT 588.530 3.670 589.070 4.280 ;
        RECT 589.910 3.670 590.450 4.280 ;
        RECT 591.290 3.670 591.830 4.280 ;
        RECT 592.670 3.670 593.210 4.280 ;
        RECT 594.050 3.670 594.590 4.280 ;
        RECT 595.430 3.670 595.970 4.280 ;
        RECT 596.810 3.670 597.350 4.280 ;
        RECT 598.190 3.670 598.730 4.280 ;
        RECT 599.570 3.670 600.110 4.280 ;
        RECT 600.950 3.670 601.490 4.280 ;
        RECT 602.330 3.670 602.870 4.280 ;
        RECT 603.710 3.670 604.250 4.280 ;
        RECT 605.090 3.670 605.630 4.280 ;
        RECT 606.470 3.670 607.010 4.280 ;
        RECT 607.850 3.670 608.390 4.280 ;
        RECT 609.230 3.670 609.770 4.280 ;
        RECT 610.610 3.670 611.150 4.280 ;
        RECT 611.990 3.670 612.530 4.280 ;
        RECT 613.370 3.670 613.910 4.280 ;
        RECT 614.750 3.670 615.290 4.280 ;
        RECT 616.130 3.670 616.670 4.280 ;
        RECT 617.510 3.670 618.050 4.280 ;
        RECT 618.890 3.670 619.430 4.280 ;
        RECT 620.270 3.670 620.810 4.280 ;
        RECT 621.650 3.670 622.190 4.280 ;
        RECT 623.030 3.670 623.570 4.280 ;
        RECT 624.410 3.670 624.950 4.280 ;
        RECT 625.790 3.670 626.330 4.280 ;
        RECT 627.170 3.670 627.710 4.280 ;
        RECT 628.550 3.670 629.090 4.280 ;
        RECT 629.930 3.670 630.470 4.280 ;
        RECT 631.310 3.670 631.850 4.280 ;
        RECT 632.690 3.670 633.230 4.280 ;
        RECT 634.070 3.670 634.610 4.280 ;
        RECT 635.450 3.670 635.990 4.280 ;
        RECT 636.830 3.670 637.370 4.280 ;
        RECT 638.210 3.670 638.750 4.280 ;
        RECT 639.590 3.670 640.130 4.280 ;
        RECT 640.970 3.670 641.510 4.280 ;
        RECT 642.350 3.670 642.890 4.280 ;
        RECT 643.730 3.670 644.270 4.280 ;
        RECT 645.110 3.670 645.650 4.280 ;
        RECT 646.490 3.670 647.030 4.280 ;
        RECT 647.870 3.670 648.410 4.280 ;
        RECT 649.250 3.670 649.790 4.280 ;
        RECT 650.630 3.670 651.170 4.280 ;
        RECT 652.010 3.670 652.550 4.280 ;
        RECT 653.390 3.670 653.930 4.280 ;
        RECT 654.770 3.670 655.310 4.280 ;
        RECT 656.150 3.670 656.690 4.280 ;
        RECT 657.530 3.670 658.070 4.280 ;
        RECT 658.910 3.670 659.450 4.280 ;
        RECT 660.290 3.670 660.830 4.280 ;
        RECT 661.670 3.670 662.210 4.280 ;
        RECT 663.050 3.670 663.590 4.280 ;
        RECT 664.430 3.670 664.970 4.280 ;
        RECT 665.810 3.670 666.350 4.280 ;
        RECT 667.190 3.670 667.730 4.280 ;
        RECT 668.570 3.670 669.110 4.280 ;
        RECT 669.950 3.670 670.490 4.280 ;
        RECT 671.330 3.670 671.870 4.280 ;
        RECT 672.710 3.670 673.250 4.280 ;
        RECT 674.090 3.670 674.630 4.280 ;
        RECT 675.470 3.670 676.010 4.280 ;
        RECT 676.850 3.670 677.390 4.280 ;
        RECT 678.230 3.670 678.770 4.280 ;
        RECT 679.610 3.670 680.150 4.280 ;
        RECT 680.990 3.670 681.530 4.280 ;
        RECT 682.370 3.670 682.910 4.280 ;
        RECT 683.750 3.670 684.290 4.280 ;
        RECT 685.130 3.670 685.670 4.280 ;
        RECT 686.510 3.670 687.050 4.280 ;
        RECT 687.890 3.670 688.430 4.280 ;
        RECT 689.270 3.670 689.810 4.280 ;
        RECT 690.650 3.670 691.190 4.280 ;
        RECT 692.030 3.670 692.570 4.280 ;
        RECT 693.410 3.670 693.950 4.280 ;
        RECT 694.790 3.670 695.330 4.280 ;
        RECT 696.170 3.670 696.710 4.280 ;
        RECT 697.550 3.670 698.090 4.280 ;
        RECT 698.930 3.670 699.470 4.280 ;
        RECT 700.310 3.670 700.850 4.280 ;
        RECT 701.690 3.670 702.230 4.280 ;
        RECT 703.070 3.670 703.610 4.280 ;
        RECT 704.450 3.670 704.990 4.280 ;
        RECT 705.830 3.670 706.370 4.280 ;
        RECT 707.210 3.670 707.750 4.280 ;
        RECT 708.590 3.670 709.130 4.280 ;
        RECT 709.970 3.670 710.510 4.280 ;
        RECT 711.350 3.670 711.890 4.280 ;
        RECT 712.730 3.670 713.270 4.280 ;
        RECT 714.110 3.670 714.650 4.280 ;
        RECT 715.490 3.670 716.030 4.280 ;
        RECT 716.870 3.670 717.410 4.280 ;
        RECT 718.250 3.670 718.790 4.280 ;
        RECT 719.630 3.670 720.170 4.280 ;
        RECT 721.010 3.670 721.550 4.280 ;
        RECT 722.390 3.670 722.930 4.280 ;
        RECT 723.770 3.670 724.310 4.280 ;
        RECT 725.150 3.670 725.690 4.280 ;
        RECT 726.530 3.670 727.070 4.280 ;
        RECT 727.910 3.670 728.450 4.280 ;
        RECT 729.290 3.670 729.830 4.280 ;
        RECT 730.670 3.670 731.210 4.280 ;
        RECT 732.050 3.670 732.590 4.280 ;
        RECT 733.430 3.670 733.970 4.280 ;
        RECT 734.810 3.670 735.350 4.280 ;
        RECT 736.190 3.670 736.730 4.280 ;
        RECT 737.570 3.670 738.110 4.280 ;
        RECT 738.950 3.670 739.490 4.280 ;
        RECT 740.330 3.670 740.870 4.280 ;
        RECT 741.710 3.670 742.250 4.280 ;
        RECT 743.090 3.670 743.630 4.280 ;
        RECT 744.470 3.670 745.010 4.280 ;
        RECT 745.850 3.670 746.390 4.280 ;
        RECT 747.230 3.670 747.770 4.280 ;
        RECT 748.610 3.670 749.150 4.280 ;
        RECT 749.990 3.670 750.530 4.280 ;
        RECT 751.370 3.670 751.910 4.280 ;
        RECT 752.750 3.670 753.290 4.280 ;
        RECT 754.130 3.670 754.670 4.280 ;
        RECT 755.510 3.670 756.050 4.280 ;
        RECT 756.890 3.670 757.430 4.280 ;
        RECT 758.270 3.670 758.810 4.280 ;
        RECT 759.650 3.670 760.190 4.280 ;
        RECT 761.030 3.670 761.570 4.280 ;
        RECT 762.410 3.670 762.950 4.280 ;
        RECT 763.790 3.670 764.330 4.280 ;
        RECT 765.170 3.670 765.710 4.280 ;
        RECT 766.550 3.670 767.090 4.280 ;
        RECT 767.930 3.670 768.470 4.280 ;
        RECT 769.310 3.670 769.850 4.280 ;
        RECT 770.690 3.670 771.230 4.280 ;
        RECT 772.070 3.670 772.610 4.280 ;
        RECT 773.450 3.670 773.990 4.280 ;
        RECT 774.830 3.670 775.370 4.280 ;
        RECT 776.210 3.670 776.750 4.280 ;
        RECT 777.590 3.670 778.130 4.280 ;
        RECT 778.970 3.670 779.510 4.280 ;
        RECT 780.350 3.670 780.890 4.280 ;
        RECT 781.730 3.670 782.270 4.280 ;
        RECT 783.110 3.670 783.650 4.280 ;
        RECT 784.490 3.670 785.030 4.280 ;
        RECT 785.870 3.670 786.410 4.280 ;
        RECT 787.250 3.670 787.790 4.280 ;
        RECT 788.630 3.670 789.170 4.280 ;
        RECT 790.010 3.670 891.570 4.280 ;
      LAYER met3 ;
        RECT 21.050 10.715 867.430 587.685 ;
  END
END counter_option1
END LIBRARY

